LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY LED7SEG IS
	GENERIC ( REFRESH_COUNTS: INTEGER := 1000 );
	PORT(	CLK: IN STD_LOGIC;
			RST: IN STD_LOGIC;
			ZEROS: IN STD_LOGIC;
			OFF: IN STD_LOGIC;
			START: IN STD_LOGIC;
			STOP: IN STD_LOGIC;
			DATA: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			SIGN: IN STD_LOGIC;------------
			DP:OUT STD_LOGIC;------------
			SEGMENTS: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			ANODES: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEH1 OF LED7SEG IS

FUNCTION F_ANODES(A: INTEGER) RETURN STD_LOGIC_VECTOR IS
VARIABLE O: STD_LOGIC_VECTOR(3 DOWNTO 0):=(OTHERS=>'1');
BEGIN
	O(A):='0';
	RETURN O;
END FUNCTION;

FUNCTION F_DIGIT4(A: STD_LOGIC_VECTOR(15 DOWNTO 0); B: INTEGER) RETURN STD_LOGIC_VECTOR IS
TYPE T_DIGITS IS ARRAY(3 DOWNTO 0) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
VARIABLE I: T_DIGITS:=(A(15 DOWNTO 12), A(11 DOWNTO 8), A(7 DOWNTO 4), A(3 DOWNTO 0));
VARIABLE O: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	O:=I(B);
	RETURN O;
END FUNCTION;

FUNCTION F_SEGMENTS(A: STD_LOGIC_VECTOR(3 DOWNTO 0)) RETURN STD_LOGIC_VECTOR IS
VARIABLE O: STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN
	CASE CONV_INTEGER(UNSIGNED(A)) IS ---G DOWNTO A
		WHEN 0 =>  O:= "1000000"; --X"3F";
		WHEN 1 =>  O:= "1111001"; --X"06";
		WHEN 2 =>  O:= "0100100"; --X"5B";
		WHEN 3 =>  O:= "0110000"; --X"4F";
		WHEN 4 =>  O:= "0011001"; --X"66";
		WHEN 5 =>  O:= "0010010"; --X"6D";
		WHEN 6 =>  O:= "0000010"; --X"7D";
		WHEN 7 =>  O:= "1111000"; --X"07";
		WHEN 8 =>  O:= "0000000"; --X"7F";
		WHEN 9 =>  O:= "0011000"; --X"67";
		WHEN 10 => O:= "0001000"; --X"77";
		WHEN 11 => O:= "0000011"; --X"7C";
		WHEN 12 => O:= "1000110"; --X"39";
		WHEN 13 => O:= "0100001"; --X"5E";
		WHEN 14 => O:= "0000110"; --X"79";
		WHEN 15 => O:= "0001110"; --X"71";
		WHEN OTHERS => O:="1111111";
	END CASE;
	RETURN O;
END FUNCTION;

SIGNAL IDX: INTEGER RANGE 0 TO 3;
SIGNAL REFRESH, KEEP_VALUE : STD_LOGIC;
SIGNAL REG_DATA, REG_DATA1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
TYPE T_STATE IS (IDLE, COUNTER);
SIGNAL STATE: T_STATE;
SIGNAL REG_DP1,REG_DP : STD_LOGIC;--------------
BEGIN
	PROCESS(CLK,RST, REFRESH)
	BEGIN
		IF RST='1' THEN
			IDX <= 3;
		ELSIF RISING_EDGE(CLK) AND REFRESH='1' THEN
			IF IDX = 0 THEN
				IDX <= 3;
			ELSE
				IDX <= IDX-1;
			END IF;
		END IF;
	END PROCESS;

	PROCESS(CLK,RST,IDX,DATA,REFRESH)
	VARIABLE DIGIT4: STD_LOGIC_VECTOR(3 DOWNTO 0);
	BEGIN
		 IF RST = '1' THEN
			 SEGMENTS <= (OTHERS=>'1');  		
			 ANODES <= (OTHERS=>'1');
			 REG_DATA1 <= (OTHERS=>'0');
			 REG_DATA <= (OTHERS=>'0');
			 KEEP_VALUE <= '0';
			 DP<='1';-------------------
		 ELSIF RISING_EDGE(CLK) AND REFRESH='1' THEN
			CASE STATE IS
				WHEN IDLE =>	
					IF OFF = '1' THEN
						ANODES<=(OTHERS=>'1');
						KEEP_VALUE <= '0';
					END IF;
					IF ZEROS = '1' THEN
						SEGMENTS <= F_SEGMENTS("0000"); 		
						ANODES <= "0000";
						KEEP_VALUE <= '0';
						DP<='1';-------------------
					END IF;	
					IF START = '1' THEN
						STATE <= COUNTER;
						KEEP_VALUE <= '0';
					END IF;
					IF KEEP_VALUE = '1' THEN
						DIGIT4 := F_DIGIT4(REG_DATA1,IDX);
						SEGMENTS <= F_SEGMENTS(DIGIT4);
						ANODES <= F_ANODES(IDX);
						DP<=REG_DP1;-------------------						
					END IF;
				WHEN OTHERS =>	
					IF OFF = '1' OR ZEROS = '1' THEN
						STATE <= IDLE;
					END IF;
					IF STOP /= '1' THEN
						REG_DATA <= DATA;			
						DIGIT4 := F_DIGIT4(REG_DATA,IDX);
						SEGMENTS <= F_SEGMENTS(DIGIT4);
						ANODES <= F_ANODES(IDX);
						REG_DP<=NOT SIGN; DP <=REG_DP;-------------------
					ELSE	
						STATE <= IDLE;
						REG_DATA1 <= REG_DATA;    	
						KEEP_VALUE <= '1';
						REG_DP1<=REG_DP;-------------------
					END IF;
			END CASE;		
		END IF;
	END PROCESS;
	
	PROCESS(CLK, RST)
		VARIABLE COUNTER: INTEGER RANGE 0 TO REFRESH_COUNTS-1;
		BEGIN
			IF RST='1' THEN
				COUNTER:= REFRESH_COUNTS-1;
				REFRESH <= '0';
			ELSIF RISING_EDGE(CLK) THEN
				IF COUNTER = 0 THEN
					COUNTER := REFRESH_COUNTS-1;
					REFRESH <= '1';
				ELSE
					COUNTER := COUNTER-1;
					REFRESH <= '0';
				END IF;
			END IF;
	END PROCESS;

END ARCHITECTURE;